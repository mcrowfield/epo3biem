configuration vga_controller_behavior_cfg of vga_controller is
   for behavior
   end for;
end vga_controller_behavior_cfg;


