configuration pos_statemachine_cfg of pos is
   for statemachine
   end for;
end pos_statemachine_cfg;


