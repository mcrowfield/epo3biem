configuration posnew_nextcopter_cfg of posnew is
   for nextcopter
   end for;
end posnew_nextcopter_cfg;


