configuration divider_behavior_cfg of divider is
   for behavior
   end for;
end divider_behavior_cfg;


