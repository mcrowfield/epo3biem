configuration helicopter_extracted_cfg of helicopter is
   for extracted
   end for;
end helicopter_extracted_cfg;


