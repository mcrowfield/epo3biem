configuration draw_renderer_cfg of draw is
   for renderer
   end for;
end draw_renderer_cfg;


